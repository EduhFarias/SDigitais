LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY LOGIC_OR IS
    PORT(
        A: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        B: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        RESULT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END LOGIC_OR;    

ARCHITECTURE EXEC OF LOGIC_OR IS
    BEGIN
        PROCESS(A, B)
        BEGIN
			RESULT <= A OR B;
        END PROCESS;
    END EXEC;
