LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ADDER IS
    PORT(
        A: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        B: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        RESULT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END ADDER;    

ARCHITECTURE EXEC OF ADDER IS
    BEGIN
        PROCESS(A, B)
        BEGIN
			RESULT <= A + B;
        END PROCESS;
    END EXEC;
