LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY REGISTERS IS
    PORT(
		C_BUS 	   :	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLK        :	IN STD_LOGIC;
		LOAD       :	IN STD_LOGIC;
		CLEAR      :	IN STD_LOGIC;
		B_BUS,A_BUS:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		CONTROLLER :    IN STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END REGISTERS;    

ARCHITECTURE EXEC OF REGISTERS IS
	 
	 SIGNAL MAR_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL MDR_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL PC_OUT : STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL MBR_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL SP_OUT : STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL LV_OUT : STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL CPP_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL TOS_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL OPC_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL H_OUT  : STD_LOGIC_VECTOR(3 DOWNTO 0);
	 
	 BEGIN
	 MAR: ENTITY WORK.MAR(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, MAR_OUT
	 );
	 
	 MDR: ENTITY WORK.MDR(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, MDR_OUT
	 );
	 
	 PC: ENTITY WORK.PC(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, PC_OUT
	 );
	 
	 MBR: ENTITY WORK.MBR(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, MBR_OUT
	 );
    
	 SP: ENTITY WORK.SP(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, SP_OUT
	 );
	 
	 LV: ENTITY WORK.LV(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, LV_OUT
	 );
	 
	 CPP: ENTITY WORK.CPP(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, CPP_OUT
	 );
	 
	 TOS: ENTITY WORK.TOS(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, TOS_OUT
	 );
	 
	 OPC: ENTITY WORK.OPC(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, OPC_OUT
	 );
	 
	 H: ENTITY WORK.H(EXEC) PORT MAP(
		C_BUS, CLK, LOAD, CLEAR, H_OUT
	 );
	 
	 --ADD UM CONTROLLER PARA SELECIONAR O REGISTRADOR 
    PROCESS(CONTROLLER)
        BEGIN
	    A_BUS <= H_OUT; -- DIRECIONA PARA ENTRADA 'A' DA ULA 
		
            CASE CONTROLLER IS
                WHEN "0000" =>
                    B_BUS <= MDR_OUT;
                WHEN "0001" =>
                    B_BUS <= PC_OUT;
                WHEN "0010" =>
                    B_BUS <= MBR_OUT;
                WHEN "0011" =>
                    B_BUS <= MBRU_OUT;
                WHEN "0100" =>
                    B_BUS <= SP_OUT;
		WHEN "0101" =>
                    B_BUS <= LV_OUT;
		WHEN "0111" =>
                    B_BUS <= CPP_OUT;
		WHEN "1000" =>
                    B_BUS <= TOS_OUT;
		WHEN "1001" =>
                    B_BUS <= OPC_OUT;	  
		WHEN OTHERS =>
                    B_BUS <= "XXXX";
            END CASE;
        END PROCESS;
    END EXEC;
