LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY SUB IS
    PORT(
        A: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        RESULT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END SUB;    

ARCHITECTURE EXEC OF SUB IS
    BEGIN
        PROCESS(A, B)
        BEGIN
			RESULT <= A + (NOT B) + 1;
        END PROCESS;
    END EXEC;