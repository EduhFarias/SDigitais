LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY REGISTERS IS
    PORT(
		DATA_INPUT :	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLK        :	IN STD_LOGIC;
		LOAD       :	IN STD_LOGIC;
		CLEAR      :	IN STD_LOGIC;
		DATA_OUTPUT:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END REGISTERS;    

ARCHITECTURE EXEC OF REGISTERS IS
	 
	 SIGNAL MAR_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL MDR_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL PC_OUT : STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL MBR_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL SP_OUT : STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL LV_OUT : STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL CPP_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL TOS_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL OPC_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL H_OUT  : STD_LOGIC_VECTOR(3 DOWNTO 0);
	 
	 BEGIN
	 MAR: ENTITY WORK.MAR(EXEC) PORT MAP(
		DATA_INPUT, CLK, LOAD, CLEAR, MAR_OUT
	 );
	 
	 MDR: ENTITY WORK.MDR(EXEC) PORT MAP(
		DATA_INPUT, CLK, LOAD, CLEAR, MDR_OUT
	 );
	 
	 PC: ENTITY WORK.PC(EXEC) PORT MAP(
		DATA_INPUT, CLK, LOAD, CLEAR, PC_OUT
	 );
	 
	 MBR: ENTITY WORK.MBR(EXEC) PORT MAP(
		DATA_INPUT, CLK, LOAD, CLEAR, MBR_OUT
	 );
    
	 SP: ENTITY WORK.SP(EXEC) PORT MAP(
		DATA_INPUT, CLK, LOAD, CLEAR, SP_OUT
	 );
	 
	 LV: ENTITY WORK.LV(EXEC) PORT MAP(
		DATA_INPUT, CLK, LOAD, CLEAR, LV_OUT
	 );
	 
	 CPP: ENTITY WORK.CPP(EXEC) PORT MAP(
		DATA_INPUT, CLK, LOAD, CLEAR, CPP_OUT
	 );
	 
	 TOS: ENTITY WORK.TOS(EXEC) PORT MAP(
		DATA_INPUT, CLK, LOAD, CLEAR, TOS_OUT
	 );
	 
	 OPC: ENTITY WORK.OPC(EXEC) PORT MAP(
		DATA_INPUT, CLK, LOAD, CLEAR, OPC_OUT
	 );
	 
	 H: ENTITY WORK.H(EXEC) PORT MAP( -- COLOCAR SAIDA NA ULA
		DATA_INPUT, CLK, LOAD, CLEAR, H_OUT
	 );
	 
	 --ADD UM CONTROLLER PARA SELECIONAR O REGISTRADOR 
    PROCESS(CONTROLLER)
        BEGIN
            CASE CONTROLLER IS
                WHEN "0000" =>
                    DATA_OUTPUT <= MAR_OUT;
                WHEN "0001" =>
                    DATA_OUTPUT <= MDR_OUT;
                WHEN "0010" =>
                    DATA_OUTPUT <= PC_OUT;
                WHEN "0011" =>
                    DATA_OUTPUT <= MBR_OUT;
                WHEN "0100" =>
                    DATA_OUTPUT <= SP_OUT;
					 WHEN "0101" =>
                    DATA_OUTPUT <= LV_OUT;
					 WHEN "0111" =>
                    DATA_OUTPUT <= CPP_OUT;
					 WHEN "1000" =>
                    DATA_OUTPUT <= TOS_OUT;
					 WHEN "1001" =>
                    DATA_OUTPUT <= OPC_OUT;
					 WHEN "1010" =>
                    DATA_OUTPUT <= H_OUT;	  
					 WHEN OTHERS =>
                    RESULT <= "XXXX";
            END CASE;
        END PROCESS;
    END EXEC;
