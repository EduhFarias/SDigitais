LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MBR IS
	PORT(
		DATA_INPUT :	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLK :	IN STD_LOGIC;
		LOAD :	IN STD_LOGIC;
		CLEAR :	IN STD_LOGIC;
		DATA_OUTPUT :	OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END MBR;

ARCHITECTURE EXEC OF REG IS

	SIGNAL MIX_OUT : STD_LOGIC_VECTOR(8 DOWNTO 0);
	
BEGIN
	
   PROCESS(DATA_INPUT, CLK, LOAD, CLEAR)
   BEGIN

		IF CLEAR = '1' THEN
					DATA_OUTPUT <= "0";
		ELSIF RISING_EDGE(CLK) THEN
			IF LOAD = '1' THEN
				MIX_OUT <= MIX_OUT(3 DOWNTO 0) & DATA_INPUT;
			END IF;
		END IF;
		DATA_OUTPUT <= DATA_OUTPUT & MIX_OUT;
   END PROCESS;
    
END EXEC;
