LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY REG IS
	port(	
		DATA_INPUT :	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLK :	IN STD_LOGIC;
		LOAD :	IN STD_LOGIC;
		CLEAR:	IN STD_LOGIC;
		DATA_OUTPUT:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END REG;


ARCHITECTURE EXEC OF REG IS

    SIGNAL DO_TEMP : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

    PROCESS(I, CLK, LOAD, CLEAR)
    BEGIN

	IF CLEAR = '0' THEN
            DO_TEMP <= (DO_TEMP'RANGE => '0');
	ELSIF (CLK = '1' AND CLK'EVENT) THEN
	    IF LOAD = '1' THEN
		DO_TEMP <= DATA_INPUT;
	    END IF;
	END IF;

    END PROCESS;
    DATA_OUTPUT <= DO_TEMP;

END EXEC;
