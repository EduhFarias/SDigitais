LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY MANAGER IS
	PORT(
		A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		B : IN STD_LOGIC_VECTOR(31 DOWNTO 0)
		
	);
END MANAGER;

ARCHITECTURE EXEC OF MANAGER IS

SIGNAL ALU_OUT 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL CONTROL_ALU: STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL REG_OUT 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL CONTROL_REG: STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN 
	ALU: ENTITY WORK.BEHV PORT MAP(A, B, CONTROL_ALU, ALU_OUT);
	REG: ENTITY WORK.EXEC PORT MAP(ALU_OUT, CONTROL_REG);
	
END EXEC;
