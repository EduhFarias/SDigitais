-- Shifter

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SHFT IS
	port(	
		CLK :	IN STD_LOGIC;
		INPUT :	IN STD_LOGIC;
		CLEAR :	IN STD_LOGIC;
		DATA_OUTPUT :	OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END SHFT;


ARCHITECTURE EXEC OF SHFT IS
SIGNAL D_OUT : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
    PROCESS(INPUT, CLK, CLEAR)
	 BEGIN
	 IF CLEAR = '1' THEN
		DATA_OUTPUT <= "0000";
	 ELSIF RISING_EDGE(CLK) THEN
		    D_OUT(3 DOWNTO 1) <= D_OUT(2 DOWNTO 0);
			 D_OUT(0) <= INPUT;
	 END IF;
	 DATA_OUTPUT <= D_OUT;
    END PROCESS;
END EXEC;
