LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ULA IS
    PORT(
        A: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        CONTROLLER: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        RESULT: OU STD_LOGIC_VECTOR(3 DOWNTO 0);
    );
END ULA;    

ARCHITECTURE EXEC OF ULA IS
    BEGIN
        PROCESS(A, B ,CONTROLLER)
        BEGIN
            CASE CONTROLLER IS
                WHEN "000" =>
                    RESULT <= A + B;
                WHEN "001" =>
                    RESULT <= A + (NOT B) + 1;
                WHEN "010" =>
                    RESULT <= A AND B;
                WHEN "011" =>
                    RESULT <= A OR B
                WHEN OTHERS =>
                    RESULT <= "XXXX"
            END CASE;
        END PROCESS;
    END EXEC;
