LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY REGISTERS IS
	PORT MAP(
		-- MAR, MDR, PC, MBR -> REGISTRADORES DE CONTROLE DE MEMORIA
		-- SP, LV, CPP, TOS, OPC, H E DESLOCADOR(SHIFT-REGISTER)
	);
END REGISTERS;
