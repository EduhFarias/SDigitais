LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ULA IS
    PORT(
        A: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        CONTROLLER: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        RESULT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END ULA;    

ARCHITECTURE EXEC OF ULA IS
	 
	 SIGNAL ADD_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL SUB_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL AND_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL OR_OUT: STD_LOGIC_VECTOR(3 DOWNTO 0);
	 
	 BEGIN
	 ADDER: ENTITY WORK.ADDER(EXEC) PORT MAP(
		A, B, ADD_OUT
	 );
	 
	 SUB: ENTITY WORK.SUB(EXEC) PORT MAP(
		A, B, SUB_OUT
	 );
	 
	 OP_AND: ENTITY WORK.LOGIC_AND(EXEC) PORT MAP(
		A, B, AND_OUT
	 );
	 
	 OP_OR: ENTITY WORK.LOGIC_OR(EXEC) PORT MAP(
		A, B, OR_OUT
	 );
    
    PROCESS(A, B ,CONTROLLER)
        BEGIN
            CASE CONTROLLER IS
                WHEN "000" =>
                    RESULT <= ADD_OUT;
                WHEN "001" =>
                    RESULT <= SUB_OUT;
                WHEN "010" =>
                    RESULT <= AND_OUT;
                WHEN "011" =>
                    RESULT <= OR_OUT;
                WHEN OTHERS =>
                    RESULT <= "XXXX";
            END CASE;
        END PROCESS;
    END EXEC;
