LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ULA IS
    PORT(
        A: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        RESULT: OU STD_LOGIC_VECTOR(3 DOWNTO 0);
    );
END ULA;    

ARCHITECTURE EXEC OF ULA IS
    BEGIN
        PROCESS(A, B ,CONTROLLER)
        	RESULT <= A OR B;
        END PROCESS;
    END EXEC;
