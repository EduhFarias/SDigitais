LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY LOGIC_AND IS
    PORT(
        A: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        B: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        RESULT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END LOGIC_AND;    

ARCHITECTURE EXEC OF LOGIC_AND IS
    BEGIN
        PROCESS(A, B)
		  BEGIN
			RESULT <= A AND B;
        END PROCESS;
    END EXEC;
